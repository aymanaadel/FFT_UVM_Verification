module FFT_sva(FFT_if.DUT fft_if);

	// Write your Assertions here...

endmodule