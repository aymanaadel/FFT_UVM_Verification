assign clk = fft_if.clk;
assign rst = fft_if.rst;
// input assigns
assign x0 = fft_if.x0;
assign x1 = fft_if.x1;
assign x2 = fft_if.x2;
assign x3 = fft_if.x3;
assign x4 = fft_if.x4;
assign x5 = fft_if.x5;
assign x6 = fft_if.x6;
assign x7 = fft_if.x7;
assign x8 = fft_if.x8;
assign x9 = fft_if.x9;
assign x10 = fft_if.x10;
assign x11 = fft_if.x11;
assign x12 = fft_if.x12;
assign x13 = fft_if.x13;
assign x14 = fft_if.x14;
assign x15 = fft_if.x15;
assign x16 = fft_if.x16;
assign x17 = fft_if.x17;
assign x18 = fft_if.x18;
assign x19 = fft_if.x19;
assign x20 = fft_if.x20;
assign x21 = fft_if.x21;
assign x22 = fft_if.x22;
assign x23 = fft_if.x23;
assign x24 = fft_if.x24;
assign x25 = fft_if.x25;
assign x26 = fft_if.x26;
assign x27 = fft_if.x27;
assign x28 = fft_if.x28;
assign x29 = fft_if.x29;
assign x30 = fft_if.x30;
assign x31 = fft_if.x31;
// output assigns
assign fft_if.Yr0 = Yr0;
assign fft_if.Yr1 = Yr1;
assign fft_if.Yr2 = Yr2;
assign fft_if.Yr3 = Yr3;
assign fft_if.Yr4 = Yr4;
assign fft_if.Yr5 = Yr5;
assign fft_if.Yr6 = Yr6;
assign fft_if.Yr7 = Yr7;
assign fft_if.Yr8 = Yr8;
assign fft_if.Yr9 = Yr9;
assign fft_if.Yr10 = Yr10;
assign fft_if.Yr11 = Yr11;
assign fft_if.Yr12 = Yr12;
assign fft_if.Yr13 = Yr13;
assign fft_if.Yr14 = Yr14;
assign fft_if.Yr15 = Yr15;
assign fft_if.Yr16 = Yr16;
assign fft_if.Yr17 = Yr17;
assign fft_if.Yr18 = Yr18;
assign fft_if.Yr19 = Yr19;
assign fft_if.Yr20 = Yr20;
assign fft_if.Yr21 = Yr21;
assign fft_if.Yr22 = Yr22;
assign fft_if.Yr23 = Yr23;
assign fft_if.Yr24 = Yr24;
assign fft_if.Yr25 = Yr25;
assign fft_if.Yr26 = Yr26;
assign fft_if.Yr27 = Yr27;
assign fft_if.Yr28 = Yr28;
assign fft_if.Yr29 = Yr29;
assign fft_if.Yr30 = Yr30;
assign fft_if.Yr31 = Yr31;
assign fft_if.Yi0 = Yi0;
assign fft_if.Yi1 = Yi1;
assign fft_if.Yi2 = Yi2;
assign fft_if.Yi3 = Yi3;
assign fft_if.Yi4 = Yi4;
assign fft_if.Yi5 = Yi5;
assign fft_if.Yi6 = Yi6;
assign fft_if.Yi7 = Yi7;
assign fft_if.Yi8 = Yi8;
assign fft_if.Yi9 = Yi9;
assign fft_if.Yi10 = Yi10;
assign fft_if.Yi11 = Yi11;
assign fft_if.Yi12 = Yi12;
assign fft_if.Yi13 = Yi13;
assign fft_if.Yi14 = Yi14;
assign fft_if.Yi15 = Yi15;
assign fft_if.Yi16 = Yi16;
assign fft_if.Yi17 = Yi17;
assign fft_if.Yi18 = Yi18;
assign fft_if.Yi19 = Yi19;
assign fft_if.Yi20 = Yi20;
assign fft_if.Yi21 = Yi21;
assign fft_if.Yi22 = Yi22;
assign fft_if.Yi23 = Yi23;
assign fft_if.Yi24 = Yi24;
assign fft_if.Yi25 = Yi25;
assign fft_if.Yi26 = Yi26;
assign fft_if.Yi27 = Yi27;
assign fft_if.Yi28 = Yi28;
assign fft_if.Yi29 = Yi29;
assign fft_if.Yi30 = Yi30;
assign fft_if.Yi31 = Yi31;
