seq_item.rst=0;
seq_item.x0=16'd256;
seq_item.x1=16'd256;
seq_item.x2=16'd256;
seq_item.x3=16'd256; 
seq_item.x4=16'd256; 
seq_item.x5=16'd256;   
seq_item.x6=16'd256; 
seq_item.x7=16'd256;
seq_item.x8=16'd256;   
seq_item.x9=16'd256; 
seq_item.x10=16'd256;  
seq_item.x11=16'd256; 
seq_item.x12=16'd256;  
seq_item.x13=16'd256; 
seq_item.x14=16'd256; 
seq_item.x15=16'd256;
seq_item.x16=16'd256;  
seq_item.x17=16'd256; 
seq_item.x18=16'd256;  
seq_item.x19=16'd256; 
seq_item.x20=16'd256; 
seq_item.x21=16'd256; 
seq_item.x22=16'd256; 
seq_item.x23=16'd256;
seq_item.x24=16'd256;  
seq_item.x25=16'd256; 
seq_item.x26 =16'd256; 
seq_item.x27 =16'd256; 
seq_item.x28 =16'd256; 
seq_item.x29 =16'd256; 
seq_item.x30 =16'd256; 
seq_item.x31=16'd256;
