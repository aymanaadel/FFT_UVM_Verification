$sformat(x_str[0], "%b", seq_item.x0);
$sformat(x_str[1], "%b", seq_item.x1);
$sformat(x_str[2], "%b", seq_item.x2);
$sformat(x_str[3], "%b", seq_item.x3);
$sformat(x_str[4], "%b", seq_item.x4);
$sformat(x_str[5], "%b", seq_item.x5);
$sformat(x_str[6], "%b", seq_item.x6);
$sformat(x_str[7], "%b", seq_item.x7);
$sformat(x_str[8], "%b", seq_item.x8);
$sformat(x_str[9], "%b", seq_item.x9);
$sformat(x_str[10], "%b", seq_item.x10);
$sformat(x_str[11], "%b", seq_item.x11);
$sformat(x_str[12], "%b", seq_item.x12);
$sformat(x_str[13], "%b", seq_item.x13);
$sformat(x_str[14], "%b", seq_item.x14);
$sformat(x_str[15], "%b", seq_item.x15);
$sformat(x_str[16], "%b", seq_item.x16);
$sformat(x_str[17], "%b", seq_item.x17);
$sformat(x_str[18], "%b", seq_item.x18);
$sformat(x_str[19], "%b", seq_item.x19);
$sformat(x_str[20], "%b", seq_item.x20);
$sformat(x_str[21], "%b", seq_item.x21);
$sformat(x_str[22], "%b", seq_item.x22);
$sformat(x_str[23], "%b", seq_item.x23);
$sformat(x_str[24], "%b", seq_item.x24);
$sformat(x_str[25], "%b", seq_item.x25);
$sformat(x_str[26], "%b", seq_item.x26);
$sformat(x_str[27], "%b", seq_item.x27);
$sformat(x_str[28], "%b", seq_item.x28);
$sformat(x_str[29], "%b", seq_item.x29);
$sformat(x_str[30], "%b", seq_item.x30);
$sformat(x_str[31], "%b", seq_item.x31);
$sformat(Yr_str[0], "%b", seq_item.Yr0);
$sformat(Yr_str[1], "%b", seq_item.Yr1);
$sformat(Yr_str[2], "%b", seq_item.Yr2);
$sformat(Yr_str[3], "%b", seq_item.Yr3);
$sformat(Yr_str[4], "%b", seq_item.Yr4);
$sformat(Yr_str[5], "%b", seq_item.Yr5);
$sformat(Yr_str[6], "%b", seq_item.Yr6);
$sformat(Yr_str[7], "%b", seq_item.Yr7);
$sformat(Yr_str[8], "%b", seq_item.Yr8);
$sformat(Yr_str[9], "%b", seq_item.Yr9);
$sformat(Yr_str[10], "%b", seq_item.Yr10);
$sformat(Yr_str[11], "%b", seq_item.Yr11);
$sformat(Yr_str[12], "%b", seq_item.Yr12);
$sformat(Yr_str[13], "%b", seq_item.Yr13);
$sformat(Yr_str[14], "%b", seq_item.Yr14);
$sformat(Yr_str[15], "%b", seq_item.Yr15);
$sformat(Yr_str[16], "%b", seq_item.Yr16);
$sformat(Yr_str[17], "%b", seq_item.Yr17);
$sformat(Yr_str[18], "%b", seq_item.Yr18);
$sformat(Yr_str[19], "%b", seq_item.Yr19);
$sformat(Yr_str[20], "%b", seq_item.Yr20);
$sformat(Yr_str[21], "%b", seq_item.Yr21);
$sformat(Yr_str[22], "%b", seq_item.Yr22);
$sformat(Yr_str[23], "%b", seq_item.Yr23);
$sformat(Yr_str[24], "%b", seq_item.Yr24);
$sformat(Yr_str[25], "%b", seq_item.Yr25);
$sformat(Yr_str[26], "%b", seq_item.Yr26);
$sformat(Yr_str[27], "%b", seq_item.Yr27);
$sformat(Yr_str[28], "%b", seq_item.Yr28);
$sformat(Yr_str[29], "%b", seq_item.Yr29);
$sformat(Yr_str[30], "%b", seq_item.Yr30);
$sformat(Yr_str[31], "%b", seq_item.Yr31);
$sformat(Yi_str[0], "%b", seq_item.Yi0);
$sformat(Yi_str[1], "%b", seq_item.Yi1);
$sformat(Yi_str[2], "%b", seq_item.Yi2);
$sformat(Yi_str[3], "%b", seq_item.Yi3);
$sformat(Yi_str[4], "%b", seq_item.Yi4);
$sformat(Yi_str[5], "%b", seq_item.Yi5);
$sformat(Yi_str[6], "%b", seq_item.Yi6);
$sformat(Yi_str[7], "%b", seq_item.Yi7);
$sformat(Yi_str[8], "%b", seq_item.Yi8);
$sformat(Yi_str[9], "%b", seq_item.Yi9);
$sformat(Yi_str[10], "%b", seq_item.Yi10);
$sformat(Yi_str[11], "%b", seq_item.Yi11);
$sformat(Yi_str[12], "%b", seq_item.Yi12);
$sformat(Yi_str[13], "%b", seq_item.Yi13);
$sformat(Yi_str[14], "%b", seq_item.Yi14);
$sformat(Yi_str[15], "%b", seq_item.Yi15);
$sformat(Yi_str[16], "%b", seq_item.Yi16);
$sformat(Yi_str[17], "%b", seq_item.Yi17);
$sformat(Yi_str[18], "%b", seq_item.Yi18);
$sformat(Yi_str[19], "%b", seq_item.Yi19);
$sformat(Yi_str[20], "%b", seq_item.Yi20);
$sformat(Yi_str[21], "%b", seq_item.Yi21);
$sformat(Yi_str[22], "%b", seq_item.Yi22);
$sformat(Yi_str[23], "%b", seq_item.Yi23);
$sformat(Yi_str[24], "%b", seq_item.Yi24);
$sformat(Yi_str[25], "%b", seq_item.Yi25);
$sformat(Yi_str[26], "%b", seq_item.Yi26);
$sformat(Yi_str[27], "%b", seq_item.Yi27);
$sformat(Yi_str[28], "%b", seq_item.Yi28);
$sformat(Yi_str[29], "%b", seq_item.Yi29);
$sformat(Yi_str[30], "%b", seq_item.Yi30);
$sformat(Yi_str[31], "%b", seq_item.Yi31);
