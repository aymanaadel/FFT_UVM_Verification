rsp_seq_item.rst=FFT_vif.rst;
// inputs
rsp_seq_item.x0=FFT_vif.x0;
rsp_seq_item.x1=FFT_vif.x1;
rsp_seq_item.x2=FFT_vif.x2;
rsp_seq_item.x3=FFT_vif.x3;
rsp_seq_item.x4=FFT_vif.x4;
rsp_seq_item.x5=FFT_vif.x5;
rsp_seq_item.x6=FFT_vif.x6;
rsp_seq_item.x7=FFT_vif.x7;
rsp_seq_item.x8=FFT_vif.x8;
rsp_seq_item.x9=FFT_vif.x9;
rsp_seq_item.x10=FFT_vif.x10;
rsp_seq_item.x11=FFT_vif.x11;
rsp_seq_item.x12=FFT_vif.x12;
rsp_seq_item.x13=FFT_vif.x13;
rsp_seq_item.x14=FFT_vif.x14;
rsp_seq_item.x15=FFT_vif.x15;
rsp_seq_item.x16=FFT_vif.x16;
rsp_seq_item.x17=FFT_vif.x17;
rsp_seq_item.x18=FFT_vif.x18;
rsp_seq_item.x19=FFT_vif.x19;
rsp_seq_item.x20=FFT_vif.x20;
rsp_seq_item.x21=FFT_vif.x21;
rsp_seq_item.x22=FFT_vif.x22;
rsp_seq_item.x23=FFT_vif.x23;
rsp_seq_item.x24=FFT_vif.x24;
rsp_seq_item.x25=FFT_vif.x25;
rsp_seq_item.x26=FFT_vif.x26;
rsp_seq_item.x27=FFT_vif.x27;
rsp_seq_item.x28=FFT_vif.x28;
rsp_seq_item.x29=FFT_vif.x29;
rsp_seq_item.x30=FFT_vif.x30;
rsp_seq_item.x31=FFT_vif.x31;
// outputs
rsp_seq_item.Yr0=FFT_vif.Yr0;
rsp_seq_item.Yr1=FFT_vif.Yr1;
rsp_seq_item.Yr2=FFT_vif.Yr2;
rsp_seq_item.Yr3=FFT_vif.Yr3;
rsp_seq_item.Yr4=FFT_vif.Yr4;
rsp_seq_item.Yr5=FFT_vif.Yr5;
rsp_seq_item.Yr6=FFT_vif.Yr6;
rsp_seq_item.Yr7=FFT_vif.Yr7;
rsp_seq_item.Yr8=FFT_vif.Yr8;
rsp_seq_item.Yr9=FFT_vif.Yr9;
rsp_seq_item.Yr10=FFT_vif.Yr10;
rsp_seq_item.Yr11=FFT_vif.Yr11;
rsp_seq_item.Yr12=FFT_vif.Yr12;
rsp_seq_item.Yr13=FFT_vif.Yr13;
rsp_seq_item.Yr14=FFT_vif.Yr14;
rsp_seq_item.Yr15=FFT_vif.Yr15;
rsp_seq_item.Yr16=FFT_vif.Yr16;
rsp_seq_item.Yr17=FFT_vif.Yr17;
rsp_seq_item.Yr18=FFT_vif.Yr18;
rsp_seq_item.Yr19=FFT_vif.Yr19;
rsp_seq_item.Yr20=FFT_vif.Yr20;
rsp_seq_item.Yr21=FFT_vif.Yr21;
rsp_seq_item.Yr22=FFT_vif.Yr22;
rsp_seq_item.Yr23=FFT_vif.Yr23;
rsp_seq_item.Yr24=FFT_vif.Yr24;
rsp_seq_item.Yr25=FFT_vif.Yr25;
rsp_seq_item.Yr26=FFT_vif.Yr26;
rsp_seq_item.Yr27=FFT_vif.Yr27;
rsp_seq_item.Yr28=FFT_vif.Yr28;
rsp_seq_item.Yr29=FFT_vif.Yr29;
rsp_seq_item.Yr30=FFT_vif.Yr30;
rsp_seq_item.Yr31=FFT_vif.Yr31;

rsp_seq_item.Yi0=FFT_vif.Yi0;
rsp_seq_item.Yi1=FFT_vif.Yi1;
rsp_seq_item.Yi2=FFT_vif.Yi2;
rsp_seq_item.Yi3=FFT_vif.Yi3;
rsp_seq_item.Yi4=FFT_vif.Yi4;
rsp_seq_item.Yi5=FFT_vif.Yi5;
rsp_seq_item.Yi6=FFT_vif.Yi6;
rsp_seq_item.Yi7=FFT_vif.Yi7;
rsp_seq_item.Yi8=FFT_vif.Yi8;
rsp_seq_item.Yi9=FFT_vif.Yi9;
rsp_seq_item.Yi10=FFT_vif.Yi10;
rsp_seq_item.Yi11=FFT_vif.Yi11;
rsp_seq_item.Yi12=FFT_vif.Yi12;
rsp_seq_item.Yi13=FFT_vif.Yi13;
rsp_seq_item.Yi14=FFT_vif.Yi14;
rsp_seq_item.Yi15=FFT_vif.Yi15;
rsp_seq_item.Yi16=FFT_vif.Yi16;
rsp_seq_item.Yi17=FFT_vif.Yi17;
rsp_seq_item.Yi18=FFT_vif.Yi18;
rsp_seq_item.Yi19=FFT_vif.Yi19;
rsp_seq_item.Yi20=FFT_vif.Yi20;
rsp_seq_item.Yi21=FFT_vif.Yi21;
rsp_seq_item.Yi22=FFT_vif.Yi22;
rsp_seq_item.Yi23=FFT_vif.Yi23;
rsp_seq_item.Yi24=FFT_vif.Yi24;
rsp_seq_item.Yi25=FFT_vif.Yi25;
rsp_seq_item.Yi26=FFT_vif.Yi26;
rsp_seq_item.Yi27=FFT_vif.Yi27;
rsp_seq_item.Yi28=FFT_vif.Yi28;
rsp_seq_item.Yi29=FFT_vif.Yi29;
rsp_seq_item.Yi30=FFT_vif.Yi30;
rsp_seq_item.Yi31=FFT_vif.Yi31;
