FFT_vif.x0=stim_seq_item.x0;
FFT_vif.x1=stim_seq_item.x1;
FFT_vif.x2=stim_seq_item.x2;
FFT_vif.x3=stim_seq_item.x3;
FFT_vif.x4=stim_seq_item.x4;
FFT_vif.x5=stim_seq_item.x5;
FFT_vif.x6=stim_seq_item.x6;
FFT_vif.x7=stim_seq_item.x7;
FFT_vif.x8=stim_seq_item.x8;
FFT_vif.x9=stim_seq_item.x9;
FFT_vif.x10=stim_seq_item.x10;
FFT_vif.x11=stim_seq_item.x11;
FFT_vif.x12=stim_seq_item.x12;
FFT_vif.x13=stim_seq_item.x13;
FFT_vif.x14=stim_seq_item.x14;
FFT_vif.x15=stim_seq_item.x15;
FFT_vif.x16=stim_seq_item.x16;
FFT_vif.x17=stim_seq_item.x17;
FFT_vif.x18=stim_seq_item.x18;
FFT_vif.x19=stim_seq_item.x19;
FFT_vif.x20=stim_seq_item.x20;
FFT_vif.x21=stim_seq_item.x21;
FFT_vif.x22=stim_seq_item.x22;
FFT_vif.x23=stim_seq_item.x23;
FFT_vif.x24=stim_seq_item.x24;
FFT_vif.x25=stim_seq_item.x25;
FFT_vif.x26=stim_seq_item.x26;
FFT_vif.x27=stim_seq_item.x27;
FFT_vif.x28=stim_seq_item.x28;
FFT_vif.x29=stim_seq_item.x29;
FFT_vif.x30=stim_seq_item.x30;
FFT_vif.x31=stim_seq_item.x31;
