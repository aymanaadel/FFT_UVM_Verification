$sformat(x_str[0], "%b", seq_item.x0);
$sformat(x_str[1], "%b", seq_item.x1);
$sformat(x_str[2], "%b", seq_item.x2);
$sformat(x_str[3], "%b", seq_item.x3);
$sformat(x_str[4], "%b", seq_item.x4);
$sformat(x_str[5], "%b", seq_item.x5);
$sformat(x_str[6], "%b", seq_item.x6);
$sformat(x_str[7], "%b", seq_item.x7);
$sformat(x_str[8], "%b", seq_item.x8);
$sformat(x_str[9], "%b", seq_item.x9);
$sformat(x_str[10], "%b", seq_item.x10);
$sformat(x_str[11], "%b", seq_item.x11);
$sformat(x_str[12], "%b", seq_item.x12);
$sformat(x_str[13], "%b", seq_item.x13);
$sformat(x_str[14], "%b", seq_item.x14);
$sformat(x_str[15], "%b", seq_item.x15);
$sformat(x_str[16], "%b", seq_item.x16);
$sformat(x_str[17], "%b", seq_item.x17);
$sformat(x_str[18], "%b", seq_item.x18);
$sformat(x_str[19], "%b", seq_item.x19);
$sformat(x_str[20], "%b", seq_item.x20);
$sformat(x_str[21], "%b", seq_item.x21);
$sformat(x_str[22], "%b", seq_item.x22);
$sformat(x_str[23], "%b", seq_item.x23);
$sformat(x_str[24], "%b", seq_item.x24);
$sformat(x_str[25], "%b", seq_item.x25);
$sformat(x_str[26], "%b", seq_item.x26);
$sformat(x_str[27], "%b", seq_item.x27);
$sformat(x_str[28], "%b", seq_item.x28);
$sformat(x_str[29], "%b", seq_item.x29);
$sformat(x_str[30], "%b", seq_item.x30);
$sformat(x_str[31], "%b", seq_item.x31);