parameter w0r=16'd256;// 1
parameter w0i=16'd0;    // 0

parameter w1r=16'd251; // 0.981
parameter w1i=-16'd50; // -0.195

parameter w2r=16'd237; // 0.924
parameter w2i=-16'd98; // 0.383

parameter w3r=16'd213; // 0.831
parameter w3i=-16'd142; // 0.556

parameter w4r=16'd181; // 0.707
parameter w4i=-16'd181; // 0.707 

parameter w5r=16'd142; // 0.556
parameter w5i=-16'd213; // 0.831

parameter w6r=16'd98; // 0.383
parameter w6i=-16'd237; // 0.924

parameter w7r=16'd50; // 0.195
parameter w7i=-16'd251; // 0.981

parameter w8r=16'd0; // 0
parameter w8i=-16'd256; // 1

parameter w9r=-16'd50; // 0.195
parameter w9i=-16'd251; // 0.981

parameter w10r=-16'd98; // 0.383
parameter w10i=-16'd237; // 0.924

parameter w11r=-16'd142; // 0.556
parameter w11i=-16'd213; // 0.831

parameter w12r=-16'd181; // 0.707
parameter w12i=-16'd181; // 0.707

parameter w13r=-16'd213; // 0.831
parameter w13i=-16'd142; // 0.556

parameter w14r=-16'd237; // 0.924
parameter w14i=-16'd98; // 0.383

parameter w15r=-16'd251; // 0.981
parameter w15i=-16'd50; // 0.195
